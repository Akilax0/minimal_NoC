module pkt_proc();




endmodule