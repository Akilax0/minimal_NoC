module ni_tb();




endmodule;