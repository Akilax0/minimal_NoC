module async_fifo (
    ports
);
    
endmodule