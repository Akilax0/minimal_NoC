module async_fifo();




endmodule


n0 = 